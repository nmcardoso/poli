--------------------------------------------------------------------------------
-- TENTATIVAS:
-- 01: #24102 (10)
--------------------------------------------------------------------------------


library IEEE;
use IEEE.numeric_bit.all;

entity rom is
  port (
    addr: in bit_vector(3 downto 0);
    data: out bit_vector(31 downto 0)
   );
end rom;

architecture rom_arch of rom is
  type mem_tipo is array (0 to 15) of bit_vector(31 downto 0);

  -- Type R: [opcode (11b), Rm (5b), shamt (6b), Rn (5b), Rd (5b)]
  -- Type D: [opcode (11b), addr (9b), op2 (2b), Rn (5b), Rt (5b)]

  -- Fibonacci Sequence Program
  -- LDUR X0, [XZR, 0]    11111000010 000000000 00 11111 00000
  -- LDUR X1, [XZR, 8]    11111000010 000001000 00 11111 00001
  -- LDUR X2, [X31, 16]   11111000010 000010000 00 11111 00010
  -- LDUR X3, [X31, 24]   11111000010 000011000 00 11111 00011
  -- ADD X5, X1, X0       10001011000 00000 000000 00001 00101
  -- ADD X0, X1, X31      10001011000 11111 000000 00001 00000
  -- ADD X1, X5, X31      10001011000 11111 000000 00101 00001
  -- SUB X2, X2, X3       11001011000 00011 000000 00010 00010
  -- CBZ X2, L1           10110100 0000000000000000010 00010
  -- B L0                 000101 11111111111111111111111011
  -- STUR X1, [X31, 32]   11111000000 000100000 00 11111 00001
  -- B L2                 000101 00000000000000000000000000

  constant mem: mem_tipo := (
    0 => "11111000010000000000001111100000", 
    1 => "11111000010000001000001111100001",
    2 => "11111000010000010000001111100010",
    3 => "11111000010000011000001111100011",
    4 => "10001011000000000000000000100101",
    5 => "10001011000111110000000000100000",
    6 => "10001011000111110000000010100001",
    7 => "11001011000000110000000001000010",
    8 => "10110100000000000000000001000010",
    9 => "00010111111111111111111111111011",
    10 => "11111000000000100000001111100001",
    11 => "00010100000000000000000000000000",
    12 => "00000000000000000000000000000000",
    13 => "00000000000000000000000000000000",
    14 => "00000000000000000000000000000000",
    15 => "00000000000000000000000000000000"
  );
begin
   data <= mem(to_integer(unsigned(addr)));
end rom_arch;
